////////////////////////////////////////////////////////////////////////////////////////////
//
//	File: BusControl.v
// Top-level file for Bus Control Logic System (LE D.1)
//
//	Created by Addison Ferrari, 21 June 2019
// Modified by J.S. Thweatt, 14 October 2019
// Modified by K.L. Cooper, 14 January 2021
// Modified by Brenden Duffy, 21 March 2021
//
//=======================================================
//  This code is generated by Terasic System Builder
//=======================================================
//
////////////////////////////////////////////////////////////////////////////////////////////////////

// DO NOT MODIFY THE MODULE AND PORT DECLARATIONs OF THIS MODULE!

module BusControl(MAX10_CLK1_50, KEY, SW, HEX0, HEX1, HEX2, HEX3, HEX4, HEX5, LEDR, DB0, DB1, DB2);
	input        MAX10_CLK1_50;									// System clock
	input  [1:0] KEY;													// DE10 Pushbuttons
	input  [9:0] SW;													// DE10 Switches 
	output [6:0] HEX0;												// DE10 Seven-segment displays
	output [6:0] HEX1;
	output [6:0] HEX2;
	output [6:0] HEX3;
	output [6:0] HEX4;
	output [6:0] HEX5;
	output [9:0] LEDR;												// DE10 LEDs
	output [7:0] DB0, DB1, DB2;									// ports added to allow debugging of val0, val1, val2 loads

// END MODULE AND PORT DECLARATION

// BEGIN WIRE DECLARATION
	
// Buttons is the output of a Finite State Machine.
// Each time that one of the DE10 pushbuttons is pressed and released, the corresponding value of BUTTONS goes high for one clock period.
//	This ensures that a single press and release of a pushbutton enables only one register transfer.
// YOU MUST USE THE VALUES FROM BUTTONS INSTEAD OF tHE VALUES FROM KEY IN YOUR IMPLEMENTATION.
	
	wire [1:0] buttons;												// DO NOT MODIFY!

// These values represent the register states.
// The synthesis keep directive will allow you to view these wires in simulation.

	wire [7:0] val0 /* synthesis keep */ ;						// DO NOT MODIFY!
	wire [7:0] val1 /* synthesis keep */ ;						// DO NOT MODIFY!
	wire [7:0] val2 /* synthesis keep */ ;						// DO NOT MODIFY!
	wire [7:0] valL /* synthesis keep */ ;						// DO NOT MODIFY!
	wire [7:0] valA /* synthesis keep */ ;						// DO NOT MODIFY!
	wire [7:0] valB /* synthesis keep */ ;						// DO NOT MODIFY!
	wire [7:0] valC /* synthesis keep */ ;						// DO NOT MODIFY!

// You MAY alter these wire declarations if you wish, or even delete them entirely.
// What you replace them with will depend on your design.

	wire [7:0] bus; 													// Input bus
	wire       load;													// Register load

// Add your other wire declarations here

	wire D0, D1, D2, D3, lD0, lD1, lD2, lD3, Dl;
	wire [7:0] saveBus, loadBus, saveD3;
	
	

// END WIRE DECLARATION
	
// BEGIN TOP-LEVEL HARDWARE MODEL //
		
// Review the hardware description for the buttonpress module in buttonpress.v.
// Use BUTTONS as the control signal for your hardware instead of KEY.
//	This ensures that a single press and release of a pushbutton enables only one register transfer.
// DO NOT ALTER THE INSTANTIATIONS OF THE buttonpress MODULES!

//                 System clock   Pushbutton  Enable
	buttonpress bp1(MAX10_CLK1_50, KEY[1],     buttons[1]);
	buttonpress bp0(MAX10_CLK1_50, KEY[0],     buttons[0]);

// These seven-segment decoders show the associated 8-bit register values in hexadecimal on two seven-segment displays
// DO NOT ALTER THE INSTANTIATIONS OF THE hexDecoder_7seg MODULES!

//                    Upper Hex Display  Lower Hex Display  Register Value
	hexDecoder_7seg h1(HEX5,              HEX4,              valA);
	hexDecoder_7seg h2(HEX3,              HEX2,              valB);
	hexDecoder_7seg h3(HEX1,              HEX0,              valC);

// This continuous assignment connects the valL to the LEDs.
// DO NOT ALTER THIS CONTINUOUS ASSIGNMENT!
	
	assign LEDR = {2'b00, valL};

// These continuous assignments connect val0, val1, and val2 to the debugging ports so that val0, val1, val2 can be 
// seen in simulation. Without these connections, the synthesis keep directive is not effective. These are not 
// necessary for your bus control cicuit to work, but will make debugging easier. Use valX in simulation, not DBX.
// DO NOT ALTER THESE CONTINUOUS ASSIGNMENTS!
	
	assign DB0 = val0;
	assign DB1 = val1;
	assign DB2 = val2;
	
// Review the hardware description for the register module in register8bit.v
// Register rL acts as both r3 and rD. It should be capable of all register transfers described in the specification.
	
// CHANGE THE LOAD CONTROL and the REGISTER INPUTS as needed by the system you are trying to implement.
// DO NOT CHANGE THE CLOCK SOURCE OR THE REGISTER OUTPUT!

//                 System clock   Load control  Register inputs  Register outputs
	register8bit r0(MAX10_CLK1_50, D0,         saveBus,             val0);
	register8bit r1(MAX10_CLK1_50, D1,         saveBus,             val1);
	register8bit r2(MAX10_CLK1_50, D2,         saveBus,             val2);
	register8bit rL(MAX10_CLK1_50, Dl,         saveD3,             valL);

	register8bit rA(MAX10_CLK1_50, lD0,         loadBus,             valA);
	register8bit rB(MAX10_CLK1_50, lD1,         loadBus,             valB);
	register8bit rC(MAX10_CLK1_50, lD2,         loadBus,             valC);
		
// Instantiate all other hardware here.
// You may also add continuous assignments here.

saveBusIn(SW[7:0], buttons[0], SW[9:8], D0, D1, D2, D3, saveBus);

assign Dl = (buttons[0] == 1'b1) ? D3 : 
					(buttons[1] == 1'b1) ? lD3: 1'b0;
assign saveD3 = (buttons[0] == 1'b1) ? saveBus :
						(buttons[1] == 1'b1) ? loadBus: 1'b0;


loadBus(SW[9:8], SW[7:6], buttons[1], lD0, lD1, lD2, lD3, val0, val1, val2, valL, loadBus);

// END TOP-LEVEL HARDWARE MODEL //

endmodule

// Write the hardware models that you instantiate into the top-level module starting here.
module loadBus(destControl, sourceControl, enable, lD0, lD1, lD2, lD3, val0, val1, val2, valL, loadBus);
input [1:0] destControl, sourceControl;
input enable;
input [7:0] val0, val1, val2, valL;
output lD0, lD1, lD2, lD3;
output [7:0] loadBus;
twoByFourDecEnable saveOut(destControl[0], destControl[1], enable, lD0, lD1, lD2, lD3);  // Chooses which register recieves by decoder
assign loadBus = (sourceControl == 2'b00) ? val0 :
						(sourceControl == 2'b01) ? val1 :
						(sourceControl == 2'b10) ? val2 :
						(sourceControl == 2'b11) ? valL: 8'b0000_0000;

endmodule

module saveBusIn(data, enable, control, D0, D1, D2, D3, saveBus);
input [7:0] data;
input [1:0] control;
input enable;
output D0, D1, D2, D3;
output [7:0] saveBus;
twoByFourDecEnable saveOut(control[0], control[1], enable, D0, D1, D2, D3);  // Chooses which register recieves by decoder
assign saveBus = data;
endmodule


module twoByFourDecEnable(A0, A1, enable, D0, D1, D2, D3);
	input A0, A1, enable; 					
	output D0, D1, D2, D3;					
	
	assign D0 = (enable)*(~A1)*(~A0);
	assign D1 = (enable)*(~A1)*(A0);
	assign D2 = (enable)*(A1)*(~A0);
	assign D3 = (enable)*(A1)*(A0);

	
	endmodule
	

